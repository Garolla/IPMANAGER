

library IEEE;
use IEEE.STD_LOGIC_1164.all;

package CONSTANTS is

constant DATA_WIDTH : integer := 16;
constant ADD_WIDTH  : integer := 6;
end CONSTANTS;

package body CONSTANTS is

 
end CONSTANTS;
